
interface system_if (input logic fast_clk, slow_clk, reset);

endinterface
