
interface tb_clk_if(input fast_clk, slow_clk);

	logic start_fast_clock;

endinterface
