
package fp;
	localparam integer WORD_LENGTH = 16;
	typedef reg [WORD_LENGTH-1:0] fpType;
	typedef reg [2*WORD_LENGTH-1:0] fpWideType;
endpackage
