
interface tb_clk_if(input fast_clk, slow_clk, reset);

	logic start_fast_clock;

endinterface
